library verilog;
use verilog.vl_types.all;
entity cryptography_vlg_vec_tst is
end cryptography_vlg_vec_tst;
