library verilog;
use verilog.vl_types.all;
entity projeto_final_logica_vlg_vec_tst is
end projeto_final_logica_vlg_vec_tst;
