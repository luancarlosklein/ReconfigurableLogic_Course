library verilog;
use verilog.vl_types.all;
entity compare_numbers_vlg_vec_tst is
end compare_numbers_vlg_vec_tst;
