library verilog;
use verilog.vl_types.all;
entity projeto_final_forca_bruta_vlg_vec_tst is
end projeto_final_forca_bruta_vlg_vec_tst;
