library verilog;
use verilog.vl_types.all;
entity sync_ram_vlg_vec_tst is
end sync_ram_vlg_vec_tst;
